atemtvs3dcpu_i : entity work.atemtvs3dcpu 
generic map (
INCLUDE_DEBUG            => INCLUDE_DEBUG, --boolean width = null
INCLUDE_MAIN_LCD         => INCLUDE_MAIN_LCD, --boolean width = null
INCLUDE_ETHSW            => INCLUDE_ETHSW, --boolean width = null
INCLUDE_PCIE             => INCLUDE_PCIE, --boolean width = null
INCLUDE_SWITCHER         => INCLUDE_SWITCHER, --boolean width = null
INCLUDE_AUD_DLY          => INCLUDE_AUD_DLY, --boolean width = null
INCLUDE_MP1              => INCLUDE_MP1, --boolean width = null
INCLUDE_MP2              => INCLUDE_MP2, --boolean width = null
INCLUDE_MC1              => INCLUDE_MC1, --boolean width = null
INCLUDE_CLOCK_DISPLAY    => INCLUDE_CLOCK_DISPLAY, --boolean width = null
INCLUDE_MV               => INCLUDE_MV, --boolean width = null
INCLUDE_AC2              => INCLUDE_AC2, --boolean width = null
INCLUDE_MCS              => INCLUDE_MCS, --boolean width = null
INCLUDE_RAM1             => INCLUDE_RAM1, --boolean width = null
INCLUDE_LCD2             => INCLUDE_LCD2, --boolean width = null
REVISION_ID              => REVISION_ID --std_logic_vector width = 8
);
port map (
fpga1_config_d0          => fpga1_config_d0, --out width = std_logic
fpga1_config_nstatus     => fpga1_config_nstatus, --in width = std_logic
fpga1_config_nconfig     => fpga1_config_nconfig, --inout width = std_logic
fpga1_config_dclk        => fpga1_config_dclk, --out width = std_logic
adbus_mclk               => adbus_mclk, --out width = std_logic
adbus_cmd                => adbus_cmd, --out width = std_logic
adbus_sclk               => adbus_sclk, --in width = std_logic
adbus_stat               => adbus_stat, --in width = std_logic
adbus_data               => adbus_data, --inout width = std_logic_vector
audio_lrck               => audio_lrck, --in width = std_logic
audio_mclk               => audio_mclk, --in width = std_logic
audio_bitclk             => audio_bitclk, --out width = std_logic
audio_refclk_fpga        => audio_refclk_fpga, --out width = std_logic
audio_power_en           => audio_power_en, --out width = std_logic
audio_rstn               => audio_rstn, --out width = std_logic
audio_rca_din            => audio_rca_din, --in width = std_logic
audio_xlr_din            => audio_xlr_din, --in width = std_logic
audio_mic_din            => audio_mic_din, --in width = std_logic
audio_control_dout       => audio_control_dout, --out width = std_logic
audio_studio_dout        => audio_studio_dout, --out width = std_logic
audio_phones_dout        => audio_phones_dout, --out width = std_logic
audio_talkback_dout      => audio_talkback_dout, --out width = std_logic
madi_in_p                => madi_in_p, --in width = std_logic
madi_in_n                => madi_in_n, --in width = std_logic
madi_out_p               => madi_out_p, --out width = std_logic
madi_out_n               => madi_out_n, --out width = std_logic
fpga_cpu_vclk_a_p        => fpga_cpu_vclk_a_p, --in width = std_logic
fpga_cpu_vclk_a_n        => fpga_cpu_vclk_a_n, --in width = std_logic
fpga_cpu_clk_100m_c_p    => fpga_cpu_clk_100m_c_p, --in width = std_logic
fpga_cpu_clk_100m_c_n    => fpga_cpu_clk_100m_c_n, --in width = std_logic
m2_a_tx_p                => m2_a_tx_p, --out width = std_logic_vector
m2_a_tx_n                => m2_a_tx_n, --out width = std_logic_vector
m2_a_rx_p                => m2_a_rx_p, --in width = std_logic_vector
m2_a_rx_n                => m2_a_rx_n, --in width = std_logic_vector
m2_b_tx_p                => m2_b_tx_p, --out width = std_logic_vector
m2_b_tx_n                => m2_b_tx_n, --out width = std_logic_vector
m2_b_rx_p                => m2_b_rx_p, --in width = std_logic_vector
m2_b_rx_n                => m2_b_rx_n, --in width = std_logic_vector
link_fc_f1_0_p           => link_fc_f1_0_p, --out width = std_logic
link_fc_f1_0_n           => link_fc_f1_0_n, --out width = std_logic
link_fc_f1_1_p           => link_fc_f1_1_p, --out width = std_logic
link_fc_f1_1_n           => link_fc_f1_1_n, --out width = std_logic
link_fc_f1_2_p           => link_fc_f1_2_p, --out width = std_logic
link_fc_f1_2_n           => link_fc_f1_2_n, --out width = std_logic
link_fc_f1_3_p           => link_fc_f1_3_p, --out width = std_logic
link_fc_f1_3_n           => link_fc_f1_3_n, --out width = std_logic
link_f1_fc_0_p           => link_f1_fc_0_p, --in width = std_logic
link_f1_fc_0_n           => link_f1_fc_0_n, --in width = std_logic
link_f1_fc_1_p           => link_f1_fc_1_p, --in width = std_logic
link_f1_fc_1_n           => link_f1_fc_1_n, --in width = std_logic
link_f1_fc_2_p           => link_f1_fc_2_p, --in width = std_logic
link_f1_fc_2_n           => link_f1_fc_2_n, --in width = std_logic
fpga_cpu_vclk_b_p        => fpga_cpu_vclk_b_p, --in width = std_logic
fpga_cpu_vclk_b_n        => fpga_cpu_vclk_b_n, --in width = std_logic
fpga_cpu_clk_100m_d_p    => fpga_cpu_clk_100m_d_p, --in width = std_logic
fpga_cpu_clk_100m_d_n    => fpga_cpu_clk_100m_d_n, --in width = std_logic
link_fc_f1_4_p           => link_fc_f1_4_p, --out width = std_logic
link_fc_f1_4_n           => link_fc_f1_4_n, --out width = std_logic
link_fc_f2_2_p           => link_fc_f2_2_p, --out width = std_logic
link_fc_f2_2_n           => link_fc_f2_2_n, --out width = std_logic
link_fc_f2_0_p           => link_fc_f2_0_p, --out width = std_logic
link_fc_f2_0_n           => link_fc_f2_0_n, --out width = std_logic
eth_int_n                => eth_int_n, --in width = std_logic
eth_rstn                 => eth_rstn, --out width = std_logic
eth_pwr_en               => eth_pwr_en, --out width = std_logic
eth_mdc                  => eth_mdc, --out width = std_logic
eth_mdio                 => eth_mdio, --inout width = std_logic
eth_clk_156m25_b_p       => eth_clk_156m25_b_p, --in width = std_logic
eth_clk_156m25_b_n       => eth_clk_156m25_b_n, --in width = std_logic
eth_usxgmiip0_txp        => eth_usxgmiip0_txp, --out width = std_logic
eth_usxgmiip0_txn        => eth_usxgmiip0_txn, --out width = std_logic
eth_usxgmiip1_txp        => eth_usxgmiip1_txp, --out width = std_logic
eth_usxgmiip1_txn        => eth_usxgmiip1_txn, --out width = std_logic
eth_usxgmiip2_txp        => eth_usxgmiip2_txp, --out width = std_logic
eth_usxgmiip2_txn        => eth_usxgmiip2_txn, --out width = std_logic
eth_usxgmiip3_txp        => eth_usxgmiip3_txp, --out width = std_logic
eth_usxgmiip3_txn        => eth_usxgmiip3_txn, --out width = std_logic
eth_usxgmiip0_rxp        => eth_usxgmiip0_rxp, --in width = std_logic
eth_usxgmiip0_rxn        => eth_usxgmiip0_rxn, --in width = std_logic
eth_usxgmiip1_rxp        => eth_usxgmiip1_rxp, --in width = std_logic
eth_usxgmiip1_rxn        => eth_usxgmiip1_rxn, --in width = std_logic
eth_usxgmiip2_rxp        => eth_usxgmiip2_rxp, --in width = std_logic
eth_usxgmiip2_rxn        => eth_usxgmiip2_rxn, --in width = std_logic
eth_usxgmiip3_rxp        => eth_usxgmiip3_rxp, --in width = std_logic
eth_usxgmiip3_rxn        => eth_usxgmiip3_rxn, --in width = std_logic
fpga_cpu_i2c_scl         => fpga_cpu_i2c_scl, --out width = std_logic
fpga_cpu_i2c_sda         => fpga_cpu_i2c_sda, --inout width = std_logic_vector
buslink_clk              => buslink_clk, --inout width = std_logic
buslink_d                => buslink_d, --inout width = std_logic_vector
auxlink_fc_f1_d          => auxlink_fc_f1_d, --inout width = std_logic_vector
auxlink_fc_f2_d          => auxlink_fc_f2_d, --inout width = std_logic_vector
fpga_cpu_clk_100m_b_p    => fpga_cpu_clk_100m_b_p, --in width = std_logic
fpga_cpu_clk_100m_b_n    => fpga_cpu_clk_100m_b_n, --in width = std_logic
fpga_cpu_ram_1_a         => fpga_cpu_ram_1_a, --out width = std_logic_vector
fpga_cpu_ram_1_act_n     => fpga_cpu_ram_1_act_n, --out width = std_logic
fpga_cpu_ram_1_ba        => fpga_cpu_ram_1_ba, --out width = std_logic_vector
fpga_cpu_ram_1_bg        => fpga_cpu_ram_1_bg, --out width = std_logic_vector
fpga_cpu_ram_1_ck_p      => fpga_cpu_ram_1_ck_p, --out width = std_logic
fpga_cpu_ram_1_ck_n      => fpga_cpu_ram_1_ck_n, --out width = std_logic
fpga_cpu_ram_1_cke       => fpga_cpu_ram_1_cke, --out width = std_logic
fpga_cpu_ram_1_cs_n      => fpga_cpu_ram_1_cs_n, --out width = std_logic
fpga_cpu_ram_1_dm        => fpga_cpu_ram_1_dm, --inout width = std_logic_vector
fpga_cpu_ram_1_odt       => fpga_cpu_ram_1_odt, --out width = std_logic
fpga_cpu_ram_1_rst_n     => fpga_cpu_ram_1_rst_n, --out width = std_logic
fpga_cpu_ram_1_dq        => fpga_cpu_ram_1_dq, --inout width = std_logic_vector
fpga_cpu_ram_1_dqs_n     => fpga_cpu_ram_1_dqs_n, --inout width = std_logic_vector
fpga_cpu_ram_1_dqs_p     => fpga_cpu_ram_1_dqs_p, --inout width = std_logic_vector
vp                       => vp, --in width = std_logic
vn                       => vn --in width = std_logic
);

atemtvs3dcpu_i : entity work.atemtvs3dcpu 
generic map (
include_debug            => include_debug, --boolean width = null
include_main_lcd         => include_main_lcd, --boolean width = null
include_ethsw            => include_ethsw, --boolean width = null
include_pcie             => include_pcie, --boolean width = null
include_switcher         => include_switcher, --boolean width = null
include_aud_dly          => include_aud_dly, --boolean width = null
include_mp1              => include_mp1, --boolean width = null
include_mp2              => include_mp2, --boolean width = null
include_mc1              => include_mc1, --boolean width = null
include_clock_display    => include_clock_display, --boolean width = null
include_mv               => include_mv, --boolean width = null
include_ac2              => include_ac2, --boolean width = null
include_mcs              => include_mcs, --boolean width = null
include_ram1             => include_ram1, --boolean width = null
include_lcd2             => include_lcd2, --boolean width = null
revision_id              => revision_id --std_logic_vector width = 8
);
port map (
clk           => clk, --in width = std_logic
probe_in0     => probe_in0, --in width = std_logic_vector
probe_out0    => probe_out0 --out width = std_logic_vector
);

